--
--  System Clock generator for ZPUINO (papilio one)
-- 
--  Copyright 2010 Alvaro Lopes <alvieboy@alvie.com>
-- 
--  Version: 1.0
-- 
--  The FreeBSD license
--  
--  Redistribution and use in source and binary forms, with or without
--  modification, are permitted provided that the following conditions
--  are met:
--  
--  1. Redistributions of source code must retain the above copyright
--     notice, this list of conditions and the following disclaimer.
--  2. Redistributions in binary form must reproduce the above
--     copyright notice, this list of conditions and the following
--     disclaimer in the documentation and/or other materials
--     provided with the distribution.
--  
--  THIS SOFTWARE IS PROVIDED BY THE AUTHOR ``AS IS'' AND ANY
--  EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
--  THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
--  PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
--  ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
--  INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
--  (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
--  OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
--  HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
--  STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
--  ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
--  ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
--

library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.VCOMPONENTS.all;

entity clkgen is
  port (
    clkin:  in std_logic;
    rstin:  in std_logic;
    clkout: out std_logic;
    clkout1: out std_logic;
    clkout2: out std_logic;
    clkvga: out  std_logic;
    clkdiv: out  std_logic;
    rstout: out std_logic
  );
end entity clkgen;

architecture behave of clkgen is

signal nclk: std_logic := '0';
signal irst: std_logic := '0';
signal vclk: std_logic := '0';

constant nclk_period: time := 10.4166666667 ns;
constant vclk_period: time := 39.583 ns;
signal divff1: std_logic := '0';
signal divff2: std_logic := '0';

begin

  nclk <= not nclk after nclk_period/2;
  vclk <= not vclk after vclk_period/2;
  clkvga <= vclk;
  clkout1 <= transport nclk after 3 ns;
  clkout <= nclk;
  rstout<=irst;
  clkdiv <= divff2;
  -- Clkdiv
  process(nclk)
  begin
    if rising_edge(nclk) then
      divff1<=not divff1;
      if divff1='1' then
        divff2<=not divff2;
      end if;
    end if;
  end process;

  process
  begin
    wait for 1 ns;
    irst<='1';
    wait until rising_edge(nclk);
    wait until rising_edge(nclk);
    wait until falling_edge(nclk);
    irst <='0';
    wait;
  end process;

end behave;
